class sequence_i extends uvm_sequence_item;

/* declaration of the item*/

    function new(string name="sequence_i",uvm_component parent=null);

        super.new(name,parent);

    endfunction

endclass