interface mem_if(input logic clk, reset);

    //define input , Define output 

    //logic 

    //logic 



endinterface